
module funcproc (
	source,
	probe);	

	output	[79:0]	source;
	input	[39:0]	probe;
endmodule
